`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:06:17 05/05/2017 
// Design Name: 
// Module Name:    encryption 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//	
//////////////////////////////////////////////////////////////////////////////////
module encryption(
		input clk,
		input [0:63] plainText,
		input [63:0] key,
		output [63:0] encrypted
    );
	
	
	reg [7:0] permInitial [63:0];
	reg [7:0] permFinal [63:0];
	reg [7:0] permExpansion [0:47];
	reg [7:0] permP [0:31];
	reg [0:3] s1 [0:3][0:15];
	reg [0:3] s2 [0:3][0:15];
	reg [0:3] s3 [0:3][0:15];
	reg [0:3] s4 [0:3][0:15];
	reg [0:3] s5 [0:3][0:15];
	reg [0:3] s6 [0:3][0:15];
	reg [0:3] s7 [0:3][0:15];
	reg [0:3] s8 [0:3][0:15];
	
	initial begin
		$readmemh("permP.data", permP);
		$readmemh("permInitial.data", permInitial);
		$readmemh("permExpansion.data", permExpansion);
		$readmemh("permFinal.data", permFinal);
	end
	
	//s1
	initial begin 
		s1[0][0]=14;
		s1[0][1]=4;
		s1[0][2]=13;
		s1[0][3]=1;
		s1[0][4]=2;
		s1[0][5]=15;
		s1[0][6]=11;
		s1[0][7]=8;
		s1[0][8]=3;
		s1[0][9]=10;
		s1[0][10]=6;
		s1[0][11]=12;
		s1[0][12]=5;
		s1[0][13]=9;
		s1[0][14]=0;
		s1[0][15]=7;
		s1[1][0]=0;
		s1[1][1]=15;
		s1[1][2]=7;
		s1[1][3]=4;
		s1[1][4]=14;
		s1[1][5]=2;
		s1[1][6]=13;
		s1[1][7]=1;
		s1[1][8]=10;
		s1[1][9]=6;
		s1[1][10]=12;
		s1[1][11]=11;
		s1[1][12]=9;
		s1[1][13]=5;
		s1[1][14]=3;
		s1[1][15]=8;
		s1[2][0]=4;
		s1[2][1]=1;
		s1[2][2]=14;
		s1[2][3]=8;
		s1[2][4]=13;
		s1[2][5]=6;
		s1[2][6]=2;
		s1[2][7]=11;
		s1[2][8]=15;
		s1[2][9]=12;
		s1[2][10]=9;
		s1[2][11]=7;
		s1[2][12]=3;
		s1[2][13]=10;
		s1[2][14]=5;
		s1[2][15]=0;
		s1[3][0]=15;
		s1[3][1]=12;
		s1[3][2]=8;
		s1[3][3]=2;
		s1[3][4]=4;
		s1[3][5]=9;
		s1[3][6]=1;
		s1[3][7]=7;
		s1[3][8]=5;
		s1[3][9]=11;
		s1[3][10]=3;
		s1[3][11]=14;
		s1[3][12]=10;
		s1[3][13]=0;
		s1[3][14]=6;
		s1[3][15]=13;
	end
	
	//s2
	initial begin
		s2[0][0]=15;
		s2[0][1]=1;
		s2[0][2]=8;
		s2[0][3]=14;
		s2[0][4]=6;
		s2[0][5]=11;
		s2[0][6]=3;
		s2[0][7]=4;
		s2[0][8]=9;
		s2[0][9]=7;
		s2[0][10]=2;
		s2[0][11]=13;
		s2[0][12]=12;
		s2[0][13]=0;
		s2[0][14]=5;
		s2[0][15]=10;
		s2[1][0]=3;
		s2[1][1]=13;
		s2[1][2]=4;
		s2[1][3]=7;
		s2[1][4]=15;
		s2[1][5]=2;
		s2[1][6]=8;
		s2[1][7]=14;
		s2[1][8]=12;
		s2[1][9]=0;
		s2[1][10]=1;
		s2[1][11]=10;
		s2[1][12]=6;
		s2[1][13]=9;
		s2[1][14]=11;
		s2[1][15]=5;
		s2[2][0]=0;
		s2[2][1]=14;
		s2[2][2]=7;
		s2[2][3]=11;
		s2[2][4]=10;
		s2[2][5]=4;
		s2[2][6]=13;
		s2[2][7]=1;
		s2[2][8]=5;
		s2[2][9]=8;
		s2[2][10]=12;
		s2[2][11]=6;
		s2[2][12]=9;
		s2[2][13]=3;
		s2[2][14]=2;
		s2[2][15]=15;
		s2[3][0]=13;
		s2[3][1]=8;
		s2[3][2]=10;
		s2[3][3]=1;
		s2[3][4]=3;
		s2[3][5]=15;
		s2[3][6]=4;
		s2[3][7]=2;
		s2[3][8]=11;
		s2[3][9]=6;
		s2[3][10]=7;
		s2[3][11]=12;
		s2[3][12]=0;
		s2[3][13]=5;
		s2[3][14]=14;
		s2[3][15]=9;
	end
	
	//s3
	initial begin
		s3[0][0]=10;
		s3[0][1]=0;
		s3[0][2]=9;
		s3[0][3]=14;
		s3[0][4]=6;
		s3[0][5]=3;
		s3[0][6]=15;
		s3[0][7]=5;
		s3[0][8]=1;
		s3[0][9]=13;
		s3[0][10]=12;
		s3[0][11]=7;
		s3[0][12]=11;
		s3[0][13]=4;
		s3[0][14]=2;
		s3[0][15]=8;
		s3[1][0]=13;
		s3[1][1]=7;
		s3[1][2]=0;
		s3[1][3]=9;
		s3[1][4]=3;
		s3[1][5]=4;
		s3[1][6]=6;
		s3[1][7]=10;
		s3[1][8]=2;
		s3[1][9]=8;
		s3[1][10]=5;
		s3[1][11]=14;
		s3[1][12]=12;
		s3[1][13]=11;
		s3[1][14]=15;
		s3[1][15]=1;
		s3[2][0]=13;
		s3[2][1]=6;
		s3[2][2]=4;
		s3[2][3]=9;
		s3[2][4]=8;
		s3[2][5]=15;
		s3[2][6]=3;
		s3[2][7]=0;
		s3[2][8]=11;
		s3[2][9]=1;
		s3[2][10]=2;
		s3[2][11]=12;
		s3[2][12]=5;
		s3[2][13]=10;
		s3[2][14]=14;
		s3[2][15]=7;
		s3[3][0]=1;
		s3[3][1]=10;
		s3[3][2]=13;
		s3[3][3]=0;
		s3[3][4]=6;
		s3[3][5]=9;
		s3[3][6]=8;
		s3[3][7]=7;
		s3[3][8]=4;
		s3[3][9]=15;
		s3[3][10]=14;
		s3[3][11]=3;
		s3[3][12]=11;
		s3[3][13]=5;
		s3[3][14]=2;
		s3[3][15]=12;
	end
	
	//s4
	initial begin
		s4[0][0]=7;
		s4[0][1]=13;
		s4[0][2]=14;
		s4[0][3]=3;
		s4[0][4]=0;
		s4[0][5]=6;
		s4[0][6]=9;
		s4[0][7]=10;
		s4[0][8]=1;
		s4[0][9]=2;
		s4[0][10]=8;
		s4[0][11]=5;
		s4[0][12]=11;
		s4[0][13]=12;
		s4[0][14]=4;
		s4[0][15]=15;
		s4[1][0]=13;
		s4[1][1]=8;
		s4[1][2]=11;
		s4[1][3]=5;
		s4[1][4]=6;
		s4[1][5]=15;
		s4[1][6]=0;
		s4[1][7]=3;
		s4[1][8]=4;
		s4[1][9]=7;
		s4[1][10]=2;
		s4[1][11]=12;
		s4[1][12]=1;
		s4[1][13]=10;
		s4[1][14]=14;
		s4[1][15]=9;
		s4[2][0]=10;
		s4[2][1]=6;
		s4[2][2]=9;
		s4[2][3]=0;
		s4[2][4]=12;
		s4[2][5]=11;
		s4[2][6]=7;
		s4[2][7]=13;
		s4[2][8]=15;
		s4[2][9]=1;
		s4[2][10]=3;
		s4[2][11]=14;
		s4[2][12]=5;
		s4[2][13]=2;
		s4[2][14]=8;
		s4[2][15]=4;
		s4[3][0]=3;
		s4[3][1]=15;
		s4[3][2]=0;
		s4[3][3]=6;
		s4[3][4]=10;
		s4[3][5]=1;
		s4[3][6]=13;
		s4[3][7]=8;
		s4[3][8]=9;
		s4[3][9]=4;
		s4[3][10]=5;
		s4[3][11]=11;
		s4[3][12]=12;
		s4[3][13]=7;
		s4[3][14]=2;
		s4[3][15]=14;
	end
	
	//s5
	initial begin
		s5[0][0]=2;
		s5[0][1]=12;
		s5[0][2]=4;
		s5[0][3]=1;
		s5[0][4]=7;
		s5[0][5]=10;
		s5[0][6]=11;
		s5[0][7]=6;
		s5[0][8]=8;
		s5[0][9]=5;
		s5[0][10]=3;
		s5[0][11]=15;
		s5[0][12]=13;
		s5[0][13]=0;
		s5[0][14]=14;
		s5[0][15]=9;
		s5[1][0]=14;
		s5[1][1]=11;
		s5[1][2]=2;
		s5[1][3]=12;
		s5[1][4]=4;
		s5[1][5]=7;
		s5[1][6]=13;
		s5[1][7]=1;
		s5[1][8]=5;
		s5[1][9]=0;
		s5[1][10]=15;
		s5[1][11]=10;
		s5[1][12]=3;
		s5[1][13]=9;
		s5[1][14]=8;
		s5[1][15]=6;
		s5[2][0]=4;
		s5[2][1]=2;
		s5[2][2]=1;
		s5[2][3]=11;
		s5[2][4]=10;
		s5[2][5]=13;
		s5[2][6]=7;
		s5[2][7]=8;
		s5[2][8]=15;
		s5[2][9]=9;
		s5[2][10]=12;
		s5[2][11]=5;
		s5[2][12]=6;
		s5[2][13]=3;
		s5[2][14]=0;
		s5[2][15]=14;
		s5[3][0]=11;
		s5[3][1]=8;
		s5[3][2]=12;
		s5[3][3]=7;
		s5[3][4]=1;
		s5[3][5]=14;
		s5[3][6]=2;
		s5[3][7]=13;
		s5[3][8]=6;
		s5[3][9]=15;
		s5[3][10]=0;
		s5[3][11]=9;
		s5[3][12]=10;
		s5[3][13]=4;
		s5[3][14]=5;
		s5[3][15]=3;
	end
	
	//s6
	initial begin
		s6[0][0]=12;
		s6[0][1]=1;
		s6[0][2]=10;
		s6[0][3]=15;
		s6[0][4]=9;
		s6[0][5]=2;
		s6[0][6]=6;
		s6[0][7]=8;
		s6[0][8]=0;
		s6[0][9]=13;
		s6[0][10]=3;
		s6[0][11]=4;
		s6[0][12]=14;
		s6[0][13]=7;
		s6[0][14]=5;
		s6[0][15]=11;
		s6[1][0]=10;
		s6[1][1]=15;
		s6[1][2]=4;
		s6[1][3]=2;
		s6[1][4]=7;
		s6[1][5]=12;
		s6[1][6]=9;
		s6[1][7]=5;
		s6[1][8]=6;
		s6[1][9]=1;
		s6[1][10]=13;
		s6[1][11]=14;
		s6[1][12]=0;
		s6[1][13]=11;
		s6[1][14]=3;
		s6[1][15]=8;
		s6[2][0]=9;
		s6[2][1]=14;
		s6[2][2]=15;
		s6[2][3]=5;
		s6[2][4]=2;
		s6[2][5]=8;
		s6[2][6]=12;
		s6[2][7]=3;
		s6[2][8]=7;
		s6[2][9]=0;
		s6[2][10]=4;
		s6[2][11]=10;
		s6[2][12]=1;
		s6[2][13]=13;
		s6[2][14]=11;
		s6[2][15]=6;
		s6[3][0]=4;
		s6[3][1]=3;
		s6[3][2]=2;
		s6[3][3]=12;
		s6[3][4]=9;
		s6[3][5]=5;
		s6[3][6]=15;
		s6[3][7]=10;
		s6[3][8]=11;
		s6[3][9]=14;
		s6[3][10]=1;
		s6[3][11]=7;
		s6[3][12]=6;
		s6[3][13]=0;
		s6[3][14]=8;
		s6[3][15]=13;
	end

	//s7
	initial begin
		s7[0][0]=4;
		s7[0][1]=11;
		s7[0][2]=2;
		s7[0][3]=14;
		s7[0][4]=15;
		s7[0][5]=0;
		s7[0][6]=8;
		s7[0][7]=13;
		s7[0][8]=3;
		s7[0][9]=12;
		s7[0][10]=9;
		s7[0][11]=7;
		s7[0][12]=5;
		s7[0][13]=10;
		s7[0][14]=6;
		s7[0][15]=1;
		s7[1][0]=13;
		s7[1][1]=0;
		s7[1][2]=11;
		s7[1][3]=7;
		s7[1][4]=4;
		s7[1][5]=9;
		s7[1][6]=1;
		s7[1][7]=10;
		s7[1][8]=14;
		s7[1][9]=3;
		s7[1][10]=5;
		s7[1][11]=12;
		s7[1][12]=2;
		s7[1][13]=15;
		s7[1][14]=8;
		s7[1][15]=6;
		s7[2][0]=1;
		s7[2][1]=4;
		s7[2][2]=11;
		s7[2][3]=13;
		s7[2][4]=12;
		s7[2][5]=3;
		s7[2][6]=7;
		s7[2][7]=14;
		s7[2][8]=10;
		s7[2][9]=15;
		s7[2][10]=6;
		s7[2][11]=8;
		s7[2][12]=0;
		s7[2][13]=5;
		s7[2][14]=9;
		s7[2][15]=2;
		s7[3][0]=6;
		s7[3][1]=11;
		s7[3][2]=13;
		s7[3][3]=8;
		s7[3][4]=1;
		s7[3][5]=4;
		s7[3][6]=10;
		s7[3][7]=7;
		s7[3][8]=9;
		s7[3][9]=5;
		s7[3][10]=0;
		s7[3][11]=15;
		s7[3][12]=14;
		s7[3][13]=2;
		s7[3][14]=3;
		s7[3][15]=12;
	end
	
	initial begin
		s8[0][0]=13;
		s8[0][1]=2;
		s8[0][2]=8;
		s8[0][3]=4;
		s8[0][4]=6;
		s8[0][5]=15;
		s8[0][6]=11;
		s8[0][7]=1;
		s8[0][8]=10;
		s8[0][9]=9;
		s8[0][10]=3;
		s8[0][11]=14;
		s8[0][12]=5;
		s8[0][13]=0;
		s8[0][14]=12;
		s8[0][15]=7;
		s8[1][0]=1;
		s8[1][1]=15;
		s8[1][2]=13;
		s8[1][3]=8;
		s8[1][4]=10;
		s8[1][5]=3;
		s8[1][6]=7;
		s8[1][7]=4;
		s8[1][8]=12;
		s8[1][9]=5;
		s8[1][10]=6;
		s8[1][11]=11;
		s8[1][12]=0;
		s8[1][13]=14;
		s8[1][14]=9;
		s8[1][15]=2;
		s8[2][0]=7;
		s8[2][1]=11;
		s8[2][2]=4;
		s8[2][3]=1;
		s8[2][4]=9;
		s8[2][5]=12;
		s8[2][6]=14;
		s8[2][7]=2;
		s8[2][8]=0;
		s8[2][9]=6;
		s8[2][10]=10;
		s8[2][11]=13;
		s8[2][12]=15;
		s8[2][13]=3;
		s8[2][14]=5;
		s8[2][15]=8;
		s8[3][0]=2;
		s8[3][1]=1;
		s8[3][2]=14;
		s8[3][3]=7;
		s8[3][4]=4;
		s8[3][5]=10;
		s8[3][6]=8;
		s8[3][7]=13;
		s8[3][8]=15;
		s8[3][9]=12;
		s8[3][10]=9;
		s8[3][11]=0;
		s8[3][12]=3;
		s8[3][13]=5;
		s8[3][14]=6;
		s8[3][15]=11;
	end

	
	//s8
	initial begin
		s7[0][0]=4;
		s7[0][1]=11;
		s7[0][2]=2;
		s7[0][3]=14;
		s7[0][4]=15;
		s7[0][5]=0;
		s7[0][6]=8;
		s7[0][7]=13;
		s7[0][8]=3;
		s7[0][9]=12;
		s7[0][10]=9;
		s7[0][11]=7;
		s7[0][12]=5;
		s7[0][13]=10;
		s7[0][14]=6;
		s7[0][15]=1;
		s7[1][0]=13;
		s7[1][1]=0;
		s7[1][2]=11;
		s7[1][3]=7;
		s7[1][4]=4;
		s7[1][5]=9;
		s7[1][6]=1;
		s7[1][7]=10;
		s7[1][8]=14;
		s7[1][9]=3;
		s7[1][10]=5;
		s7[1][11]=12;
		s7[1][12]=2;
		s7[1][13]=15;
		s7[1][14]=8;
		s7[1][15]=6;
		s7[2][0]=1;
		s7[2][1]=4;
		s7[2][2]=11;
		s7[2][3]=13;
		s7[2][4]=12;
		s7[2][5]=3;
		s7[2][6]=7;
		s7[2][7]=14;
		s7[2][8]=10;
		s7[2][9]=15;
		s7[2][10]=6;
		s7[2][11]=8;
		s7[2][12]=0;
		s7[2][13]=5;
		s7[2][14]=9;
		s7[2][15]=2;
		s7[3][0]=6;
		s7[3][1]=11;
		s7[3][2]=13;
		s7[3][3]=8;
		s7[3][4]=1;
		s7[3][5]=4;
		s7[3][6]=10;
		s7[3][7]=7;
		s7[3][8]=9;
		s7[3][9]=5;
		s7[3][10]=0;
		s7[3][11]=15;
		s7[3][12]=14;
		s7[3][13]=2;
		s7[3][14]=3;
		s7[3][15]=12;
	end
	
	
	wire [47:0] sub_key1;
	wire [47:0] sub_key2;
	wire [47:0] sub_key3;
	wire [47:0] sub_key4;
	wire [47:0] sub_key5;
	wire [47:0] sub_key6;
	wire [47:0] sub_key7;
	wire [47:0] sub_key8;
	wire [47:0] sub_key9;
	wire [47:0] sub_key10;
	wire [47:0] sub_key11;
	wire [47:0] sub_key12;
	wire [47:0] sub_key13;
	wire [47:0] sub_key14;
	wire [47:0] sub_key15;
	wire [47:0] sub_key16;
	
	generateSubkeys subKeyGenerator (
    .key(key), 
    .sub_key1(sub_key1), 
    .sub_key2(sub_key2), 
    .sub_key3(sub_key3), 
    .sub_key4(sub_key4), 
    .sub_key5(sub_key5), 
    .sub_key6(sub_key6), 
    .sub_key7(sub_key7), 
    .sub_key8(sub_key8), 
    .sub_key9(sub_key9), 
    .sub_key10(sub_key10), 
    .sub_key11(sub_key11), 
    .sub_key12(sub_key12), 
    .sub_key13(sub_key13), 
    .sub_key14(sub_key14), 
    .sub_key15(sub_key15), 
    .sub_key16(sub_key16)
    );
	
	//initial permutation of plaintex
	reg [0:63] permuted_plain;
	integer i;
	
	always @(*) begin
	
		for (i = 0; i < 64; i = i + 1) begin
			permuted_plain[i] = plainText[permInitial[i] - 1'h1];
		end
	end
	
	reg [0:31] L [16:0];
	reg [0:31] R [16:0];
	reg [0:47] e [15:0];
	
	integer h, j, k, f, l, m;
	reg [0:47] xor_e [15:0];
	wire [0:47] keys_array [0:15];
	
	assign keys_array[0] = sub_key1;
	assign keys_array[1] = sub_key2;
	assign keys_array[2] = sub_key3;
	assign keys_array[3] = sub_key4;
	assign keys_array[4] = sub_key5;
	assign keys_array[5] = sub_key6;
	assign keys_array[6] = sub_key7;
	assign keys_array[7] = sub_key8;
	assign keys_array[8] = sub_key9;
	assign keys_array[9] = sub_key10;
	assign keys_array[10] = sub_key11;
	assign keys_array[11] = sub_key12;
	assign keys_array[12] = sub_key13;
	assign keys_array[13] = sub_key14;
	assign keys_array[14] = sub_key15;
	assign keys_array[15] = sub_key16;

	reg [0:5] b [0:15][0:7];
	reg [0:31] after_s_box [0:15];
	
	reg [0:1] i_dim;
	reg [0:3] j_dim;
	reg [0:31] x [0:15];
	always @(*) begin
		L[0] = permuted_plain[0:31];
		R[0] = permuted_plain[32:63];
		for (h = 0; h < 16; h = h + 1)begin
		//key expansion
			for (j = 0; j < 48; j = j + 1)begin
				e[h][j] = R[h][permExpansion[j] - 1'h1];
			end
	
		//xors
			for (k = 0; k < 48; k = k + 1)begin
				xor_e[h][k] = keys_array[h][k] ^ e[h][k];
			end
		
			for( f = 0; f < 8; f = f + 1 ) begin
				//divide xor
				{b[h][0],b[h][1],b[h][2],b[h][3],b[h][4],b[h][5],b[h][6],b[h][7]} = {xor_e[h][0:5], xor_e[h][6:11], xor_e[h][12:17], xor_e[h][18:23], xor_e[h][24:29], xor_e[h][30:35], xor_e[h][36:41],xor_e[h][42:47]};
				
				//sboxes
				/*
				m = b[h][0]*2 + b[h][5];
				n = b[h][1]*8 + b[2]*4 + b[h][3] * 2 + b[h][4];
				*/
				
			end
			/*
			{b[h][6], b[h][1]}
			b[h][1:5]*/
			after_s_box[h] = {
			s1[{b[h][0][0], b[h][0][5]}][b[h][0][1:4]],
			s2[{b[h][1][0], b[h][1][5]}][b[h][1][1:4]],
			s3[{b[h][2][0], b[h][2][5]}][b[h][2][1:4]],
			s4[{b[h][3][0], b[h][3][5]}][b[h][3][1:4]],
			s5[{b[h][4][0], b[h][4][5]}][b[h][4][1:4]],
			s6[{b[h][5][0], b[h][5][5]}][b[h][5][1:4]],
			s7[{b[h][6][0], b[h][6][5]}][b[h][6][1:4]],
			s8[{b[h][7][0], b[h][7][5]}][b[h][7][1:4]]
			};
			
			for (l = 0; l < 32; l = l + 1)begin
				x[h][l] = after_s_box[h][permP[l] - 1'h1];
			end
			for (m = 0; m < 32; m = m + 1)begin
				R[h+1][m] = x[h][m] ^ L[h][m];
			end 
			L[h+1] = R[h];
					
			

		end
		
		
	end
	
	
	
endmodule
